----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 02/24/2021 11:20:22 AM
-- Design Name: 
-- Module Name: MPG - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity MPG is
    Port ( clk : in STD_LOGIC;
           btn : in STD_LOGIC;
           enable : out STD_LOGIC);
end MPG;
architecture Behavioral of MPG is
signal Q1,Q2,Q3: STD_LOGIC := '0';
signal count : STD_LOGIC_VECTOR (1 downto 0):="00" ;
begin
    
    process (clk)
    begin
    if rising_edge(clk) then
        count <= count + 1;
    end if;    
    end process;
    
    process(clk, btn)
    begin
        if rising_edge(clk) then
            if count = x"FFFF" then
                Q1 <= btn;
            end if;
        end if;
    end process;
    
    process (clk)
    begin
    Q2 <= Q1;
    Q3 <= Q2;
    end process;   
    
    enable <= Q2 and (not Q3);
    
  

end Behavioral;
